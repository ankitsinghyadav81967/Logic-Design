`define COUNTER_UP
